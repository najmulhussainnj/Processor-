`define EXTEST 'h00
`define IDCODE	'h01
`define SAMPLE_PRELOAD 'h02
`define SCANMODE_TE 'h03
`define SCAN1 'h04
`define SCAN2 'h05
`define SCAN3 'h06
`define SCAN4 'h07
`define SCAN5 'h08
`define SCANALL 'h12
`define SCANEN 'h13
`define FULLSCANEN 'h14
`define DEBUG	'h0A
`define MBIST	'h09
`define BYPASS 'h1f
`define DTMCONTROL 'h10
`define DMIACCESS 'h11
//`define IDCODEVALUE 32'h10e31913
`define IDCODEVALUE 32'h100039D3
