`define ABSTRACTDATASTART	  'h04
`define ABSTRACTDATAEND		  'h0f
`define DMCONTROL				    'h10
`define DMSTATUS				    'h11
`define HARTINFO				    'h12
`define ABSTRACTCNTRL	      'h16
`define ABSTRACTCMD	        'h17
`define ABSTRACTCMDAUTO	    'h18
`define CONFIGSTRINGADDR0   'h19
`define CONFIGSTRINGADDR1   'h1a
`define CONFIGSTRINGADDR2   'h1b
`define CONFIGSTRINGADDR3   'h1c
`define PBSTART				      'h20
`define PBEND					      'h2f
`define AUTHENDATA			    'h30
`define SERIALCONTROL		    'h34
`define SERIALTX            'h35
`define SERIALRX            'h36
`define BUSCONTROL			    'h38
`define BUSADDRESS0			    'h39
`define BUSADDRESS1			    'h3a
`define BUSDATA0				    'h3c
`define BUSDATA1				    'h3d
