	`define Reg_width_vme	32 
	`define Reg_width_vme_slave	32 	
